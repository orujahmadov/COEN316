-- Ibstruction cache
library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity icache is
port(
  address : in std_logic_vector(4 downto 0);
  data : out std_logic_vector(31 downto 0));
end icache;

architecture ICImplementation of icache is
  type mem is array ( 0 to 31) of std_logic_vector(31 downto 0);
  constant my_rom : mem := (
    0  => "00000000010001000100000000100000",
    1  => "00000000010001000100000000100000",
    2  => "00000000010000010001000000100000",
    3  => "00000000010001000100000000100000", 
    4  => "00000000010001000100000000100000",
    5  => "00100000000000010000000000000001",
    6  => "00000000010000010001000000100000",
    7  => "00000000010001000100000000100000",
    8  => "00000000010001000100000000100000",
    9  => "00000000010001000100000000100000",
    10 => "00000000010001000100000000100000",
    11 => "00000000010001000100000000100000",
    12 => "00000000010001000100000000100000",
    13 => "00000000010001000100000000100000",
    14 => "00000000010001000100000000100000",
    15 => "00000000000000000000000000000000",
    16 => "00000000000000000000000000000000",
    17 => "00000000000000000000000000000000",
    18 => "00000000000000000000000000000000",
    19 => "00000000000000000000000000000000",
    20 => "00000000000000000000000000000000",
    21 => "00000000000000000000000000000000",
    22 => "00000000000000000000000000000000",
    23 => "00000000000000000000000000000000",
    24 => "00000000000000000000000000000000",
    25 => "00000000000000000000000000000000",
    26 => "00000000000000000000000000000000",
    27 => "00000000000000000000000000000000",
    28 => "00000000000000000000000000000000",
    29 => "00000000000000000000000000000000",
    30 => "00000000000000000000000000000000",
    31 => "11111111111111111111111111111111");

begin
   process (address)
   begin
     data <= my_rom(to_integer(unsigned(address)));
  end process;
end architecture ICImplementation;
